module hello (
    input wire A,
    output wire B
);

    // Assign A to B
    assign B = A;
    
endmodule